`timescale 1ns / 1ps

module Encoder(
    );


endmodule
