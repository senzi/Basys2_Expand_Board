`timescale 1ns / 1ps

module flashled_555(
    );


endmodule
