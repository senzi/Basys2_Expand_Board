`timescale 1ns / 1ps

module vibration(clk,rst,up,down);
input        up,down;
input        clk,rst;  


endmodule

